* D:\_Study\CSE\CSE-209\Experiment4\Figure5\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Thu Mar 27 21:34:17 2025



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
