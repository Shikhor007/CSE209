* D:\_Study\CSE\CSE-209\Experiment4\Figure9\Schematic4.sch

* Schematics Version 9.1 - Web Update 1
* Thu Mar 27 21:58:35 2025



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic4.net"
.INC "Schematic4.als"


.probe


.END
