* D:\_Study\CSE\CSE-209\Experiment4\Figure7\Schematic3.sch

* Schematics Version 9.1 - Web Update 1
* Thu Mar 27 21:48:42 2025



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic3.net"
.INC "Schematic3.als"


.probe


.END
